`timescale 1ns/1ns

// testbench
module tb();

reg CLK, RESET, EN, OPSEL;
reg [5:0] IADDR;
reg [5:0] WADDR;
reg [5:0] OADDR;
wire [5:0] STATE;
reg [511 : 0] input_data;
reg wen, ren, cen;
reg [5 : 0] addr;
wire [511 : 0] data;


systolic_array array(
	.CLK(CLK),
	.RESET(RESET),
	.EN(EN),
	.OPSEL(OPSEL),
	.IADDR(IADDR),
	.WADDR(WADDR),
	.OADDR(OADDR),
	.STATE(STATE),
	.input_data(input_data),
	.output_buffer_wen(wen),
	.output_buffer_ren(ren),
	.output_buffer_cen(cen),
	.output_buffer_addr(addr),
	.output_buffer_data(data)
	);

initial begin
        RESET = 0;
        CLK = 1;
        EN = 0;
        OPSEL = 1;
        #100 RESET = 1;
        EN = 1;
        IADDR = 32;
        WADDR = 0;
        OADDR = 0;
        wen = 1;
        ren = 0;
        cen = 1;
        addr = 0;
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        //D = 16'b0010010000000010;
        #200
        input_data = 512'h00000000_00000000_3FE66666_00000000_00000000_00000000_BF999999_00000000_00000000_00000000_00000000_00000000_00000000_C0A99999_00000000_00000000;        
        #100
        input_data = 512'h40400000_00000000_00000000_00000000_418B3333_00000000_00000000_00000000_00000000_00000000_C0A99999_00000000_00000000_00000000_00000000_BF199999;
        #100
        input_data = 512'h00000000_00000000_00000000_BF199999_00000000_00000000_00000000_00000000_40E99999_00000000_00000000_00000000_40400000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_401AC083_00000000_00000000_C0E00000_C0A99999_00000000_00000000_00000000_00000000_00000000_410CCCCC_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_BFD99999_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_BF999999_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_BFD99999_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_BF999999_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_BFD99999_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_BF999999_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_BFD99999_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_BF999999_00000000_00000000_00000000_00000000_00000000_00000000;//
        #100
        input_data = 512'h00000000_BFD99999_00000000_00000000_00000000_00000000_00000000_00000000_00000000_3F800000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_3FE66666_00000000_00000000_00000000_BF999999_00000000_00000000_00000000_00000000_BFD99999_00000000_C0A99999_00000000_00000000;        
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_BF199999_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_BFD99999_00000000_00000000_00000000_00000000_BF999999_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_C054DD2F_00000000_00000000_00000000_00000000_406CCCCC_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_BF999999_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_BFD99999_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_BFD99999_00000000_00000000_401AC083_00000000_00000000_00000000_00000000_3F800000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_418B3333_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_3F800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_406CCCCC_00000000_00000000_00000000_00000000_00000000_00000000_00000000_BFD99999_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_BF999999_00000000_00000000_00000000_C054DD2F_00000000_00000000_00000000_00000000_00000000_BFD99999_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_C1466666_00000000_00000000_00000000_00000000_00000000_00000000_00000000_406CCCCC_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_BFD99999_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_BF999999_00000000_00000000_00000000_00000000_00000000;
        #100
        input_data = 512'h00000000_00000000_00000000_BFD99999_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        
        
        
        
        
        
        
        //datain = 77;
    end

    always #50 CLK = ~CLK;

endmodule
